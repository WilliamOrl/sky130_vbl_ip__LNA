** sch_path: /home/william/projects/sky130_vbl_ip__LNA/xschem/techsweep_pfet_g5v0d10v5.sch
**.subckt techsweep_pfet_g5v0d10v5
vg GND g DC 2.5 AC 1
vd GND d 2.5
vb GND b 0
Hn GND n vd 1
XM1 d g GND b sky130_fd_pr__pfet_g5v0d10v5 L={lx} W={wx} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code


.param wx=5 lx=0.5
.noise v(n) vg lin 100 0.1 100k 100

.control
option numdgt = 3
set wr_singlescale
set wr_vecnames

compose l_vec  values 0.5 0.51 0.52 0.53 0.54
+ 0.55 0.6 0.7 0.8 0.9 1 2 3
compose vg_vec start= 0 stop=5  step=50m
compose vd_vec start= 0 stop=5  step=50m
compose vb_vec start= 0 stop=-0.4 step=-0.2

foreach var1 $&l_vec
  alterparam lx=$var1
  reset
  foreach var2 $&vg_vec
    alter vg $var2
    foreach var3 $&vd_vec
      alter vd $var3
      foreach var4 $&vb_vec
        alter vb $var4
        run
        wrdata techsweep_pfet_g5v0d10v5.txt noise1.all
        destroy all
        set appendwrite
        unset set wr_vecnames
      end
    end
  end
end
unset appendwrite

alterparam lx=0.5
reset
op
show
write techsweep_pfet_g5v0d10v5.raw
.endc


.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt


.save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[capbd]
.save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[capbs]
.save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[cdd]
.save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[cgb]
.save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[cgd]
.save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[cgg]
.save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[cgs]
.save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[css]
.save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[gds]
.save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[gm]
.save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[gmbs]
.save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[id]
.save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[l]
.save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[vbs]
.save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[vds]
.save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[vgs]
.save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[vth]
.save onoise.m.xm1.msky130_fd_pr__pfet_g5v0d10v5.id
.save onoise.m.xm1.msky130_fd_pr__pfet_g5v0d10v5.1overf
.save g d b n


**** end user architecture code
**.ends
.GLOBAL GND
.end
